magic
tech sky130A
magscale 1 2
timestamp 1729050201
<< checkpaint >>
rect -1050 -2672 1892 486
<< error_s >>
rect 23 -877 81 -871
rect 23 -911 35 -877
rect 23 -917 81 -911
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1728978904
transform 1 0 52 0 1 -1049
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1728978904
transform 1 0 421 0 1 -1093
box -211 -319 211 319
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 in
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 gnd
port 3 nsew
<< end >>
